/*
 * Module name: CSR.sv
 * Engineer: Tommy Yee
 * Description: Interrupt enable and exception status register.
 * Dependency:
 * Status: developing
 */
module CSR(
	input  logic [7:0] addr_in,
	input  logic 
	
	
	output logic       int_en,
	output logic [5:0] ex_code
);

endmodule