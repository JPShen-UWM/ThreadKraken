module MMU(
    
);


endmodule