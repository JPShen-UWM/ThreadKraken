module alu();

int a;
assign a = 5;

endmodule