/*
 * Module name: mem_cntrl
 * Engineer:
 * Description:
 * Dependency:
 * Status: developing/testing/done
 */